`ifndef GUARD_GLOBALS
`define GUARD_GLOBALS

`define P0 8'h00
`define P1 8'h11
`define P2 8'h22
`define P3 8'h33

int error = 0;   //Global Error Counter
int num_of_pkts = 5;

`endif
